LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_arith.ALL;
USE IEEE.std_logic_unsigned.ALL;
USE IEEE.numeric_std.ALL;

ENTITY ALU IS
	PORT(
		DA : IN STD_LOGIC_VECTOR (31 DOWNTO 0); -- input1
		DB : IN STD_LOGIC_VECTOR (31 DOWNTO 0); -- input2
		ALUctrl : IN STD_LOGIC_VECTOR (2 DOWNTO 0); -- function: 0 ADD, 1 SUB, 2 AND, 3 OR and 4 LI
		Dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END ALU;

ARCHITECTURE ALU_behavior OF ALU IS
	CONSTANT ADD_CTRL : STD_LOGIC_VECTOR := "000";
	CONSTANT SUB_CTRL : STD_LOGIC_VECTOR := "001";
	CONSTANT AND_CTRL : STD_LOGIC_VECTOR := "010";
	CONSTANT OR_CTRL : STD_LOGIC_VECTOR := "011";
	CONSTANT LI_CTRL : STD_LOGIC_VECTOR := "100";
	CONSTANT JMP_CTRL : STD_LOGIC_VECTOR := "101";
	CONSTANT TLBWRITE_CTRL : STD_LOGIC_VECTOR := "110";

	SIGNAL Dout_internal : STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN
Dout_internal <= DA + DB WHEN ALUctrl = ADD_CTRL
		ELSE DA - DB WHEN ALUctrl = SUB_CTRL
		ELSE DA AND DB WHEN ALUctrl = AND_CTRL
		ELSE DA OR DB WHEN ALUctrl = OR_CTRL
		ELSE DB WHEN ALUctrl = LI_CTRL
		ELSE DA + (DB(29 DOWNTO 0) & "00") WHEN ALUctrl = JMP_CTRL
		ELSE DA WHEN ALUctrl = TLBWRITE_CTRL
		ELSE "00000000000000000000000000000000";

Dout <= Dout_internal;

END ALU_behavior;
